// SPDX-FileCopyrightText: lowRISC contributors
// SPDX-License-Identifier: Apache-2.0
// SPDX-FileContributor: Hugo McNally

package pinmux_pkg;
  parameter int unsigned COMMON_PARAMETER = 3;
  parameter int unsigned DARJEELING_SPECIFIC_PARAMETER = 4;
endpackage : pinmux_pkg
