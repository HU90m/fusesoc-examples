// SPDX-FileCopyrightText: lowRISC contributors
// SPDX-License-Identifier: Apache-2.0
// SPDX-FileContributor: Hugo McNally

module top_earlgrey;
  import pinmux_pkg::EARLGREY_SPECIFIC_PARAMETER;
endmodule : top_earlgrey
