// SPDX-FileCopyrightText: lowRISC contributors
// SPDX-License-Identifier: Apache-2.0
// SPDX-FileContributor: Hugo McNally

module top_darjeeling;
  import pinmux_pkg::DARJEELING_SPECIFIC_PARAMETER;
endmodule : top_darjeeling
